`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// NAME: EDIGA SUSEELA
// Create Date: 01.08.2023 
// Module Name: half_adder_s
// 
//////////////////////////////////////////////////////////////////////////////////


module half_adder_s(
input a,b, 
output sum,carry);
xor x1(sum,a,b); 
and a1(carry,a,b); 
endmodule

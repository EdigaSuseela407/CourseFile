`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: Alu_tb
//////////////////////////////////////////////////////////////////////////////////
module Alu_tb();
reg [3:0]a,b,s;
wire [3:0]y;
Alu uut(a,b,s,y);
integer i; 
initial
begin
a<=4'b1011;//11
b<=4'b0001;//3
for(i=0;i<16;i=i+1)
begin
	s=i;
	#10;
end
end
endmodule
